library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;


entity grass_block is
port(
	h_timer		: in unsigned (0 to 4);
	v_timer		: in unsigned (0 to 4);
	R_grass		: out std_logic_vector (0 to 3);
	G_grass		: out std_logic_vector (0 to 3);
	B_grass		: out std_logic_vector (0 to 3)
--	RGB_out		: out std_logic_vector (0 to 11)
);
end grass_block;

architecture behaviour of grass_block is
type rom_type is array (0 to 959) of std_logic_vector (0 to 11);

signal sel	: std_logic_vector (0 to 9);
signal RGB	: std_logic_vector (0 to 11);
signal rom :
rom_type:=(
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001101100100",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"001001000011",
"000100110010",
"001101100100",
"001101100100",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"000100110010",
"010010000101",
"001101100100",
"000100110010",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"001101100100",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"001101100100",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001101100100",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"001101100100",
"001101100100",
"001001000011",
"000100110010",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001001000011",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"001101100100",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"001101100100",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001101100100",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"000100110010",
"001101100100",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"010010000101",
"001001000011",
"000100110010",
"010010000101",
"001001000011",
"001001000011",
"001101100100",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001101100100",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"001101100100",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"010010000101",
"001001000011",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"001101100100",
"001101100100",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001101100100",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"001101100100",
"001101100100",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"010010000101",
"001101100100",
"000100110010",
"000100110010",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001101100100",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"010010000101",
"001101100100",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"000100110010",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"000100110010",
"001001000011",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"000100110010",
"001101100100",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001101100100",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001101100100",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"010010000101",
"010010000101",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"010010000101",
"010010000101",
"000100110010",
"000100110010",
"001001000011",
"001001000011",
"010010000101",
"001101100100",
"001001000011",
"000100110010",
"000100110010",
"010010000101",
"010010000101"
);

--select correct color for pixel address
begin
	sel <= std_logic_vector(v_timer & h_timer);
	RGB <= rom(conv_integer(sel));

	R_grass(0) <= RGB(8);
	R_grass(1) <= RGB(9);
	R_grass(2) <= RGB(10);
	R_grass(3) <= RGB(11);

	G_grass(0) <= RGB(4);
	G_grass(1) <= RGB(5);
	G_grass(2) <= RGB(6);
	G_grass(3) <= RGB(7);

	B_grass(0) <= RGB(0);
	B_grass(1) <= RGB(1);
	B_grass(2) <= RGB(2);
	B_grass(3) <= RGB(3);
end behaviour;


